/*Módulo responsável pelo Fetch de instruções*/

module Pc(addr, pc_out);

input [31:0] addr;
output [31:0] pc_out;




endmodule