module InstructionMemory(
	input Clk, 
	input [31:0] Addr,
	input [15:0] Input,
	output [31:0] InstrOut
);

reg [31:0] mem [15:0];
integer clk_single_count = 0;

always @(posedge Clk) begin
	if(clk_single_count == 0) begin
		
		//*****************--FIBONACCI WITH INPUT--*****************
		mem[0] = {16'b0000010000000001, Input[15:0]};      // ADDi: $1 = $0 + Immediate Input
		mem[1] = 32'b10000000001000010000000000000000;  	// SW: $t1, 0($a1)
		//           100000_00001_00001_0000000000000000
		mem[2] = 32'b01111100001000100000000000000000;  	// LW: $t2, 0($a1)
		//           011111_00001_00010_0000000000000000
		mem[3] = 32'b00000100000000000000000000000000;     // ADDi: $t0 = $t0 + 0 //Guarda o valor 0($zero)
		//           000001_00000_00011_0000000000000000
		mem[4] = 32'b00000100000000110000000000000000;  	// ADDi: $t3 = $t0 + 0 //Guada o F0 = 0
		//           000001_00000_00100_0000000000000001
		mem[5] = 32'b00000100000001000000000000000001;  	// ADDi: $t4 = $t0 + 1 //Guarda o F1 = 1
		//           000000_00000_00010_00101_00000000000
		mem[6] = 32'b00000000000000100010100000000000; 		// ADD: $t5 = $t0 + $t2(Input)
		//           010100_00101_00000_000000000000xxxx
		mem[7] = 32'b01010000101000000000000000001101;  	// BEQ: $t5 == $t0 -> mem[13] --> LOOP Control
		//           000000_00011_00100_00110_00000000000;
		mem[8] = 32'b00000000011001000011000000000000;     // ADD: $t6 = $t3 + $t4
		//				  100001_00100_00000_0000000000000000
		mem[9] = 32'b10000100011000000000000000000000;    // PRINT: $t3
		//				 000000_00100_00000_00011_00000000000
		mem[10] = 32'b00000000100000000001100000000000;    // ADD: $t3 = $t4 + $t0
		//				  000000_00110_00000_00100_00000000000
		mem[11] = 32'b00000000110000000010000000000000;    // ADD: $t4 = $t6 + $t0
		//				  000011_00101_00101_0000000000000001;
		mem[12] = 32'b00001100101001010000000000000001;    // SUB: $t5 = $t5 - 1
		//				  010001_00000000000000000000000011
		mem[13] = 32'b010001_00000000000000000000000111;    // JUMP: Addr == 7		
		//				  100001_00100_00000_0000000000000000
		mem[14] = 32'b100001_00011_000000000000000000000;   // PRINT: $t3
		
		clk_single_count = 1;
	end
end
assign InstrOut = mem[Addr];
endmodule


		//*****************--JAL TEST--******************
		//           000001_00000_00001_0000000000000101
		//mem[0] = 32'b00000100000000010000000000000101; //ADDi: $1 = $0 + 5
		//           000001_00000_00010_0000000000001010
		//mem[1] = 32'b00000100000000100000000000001010; //ADDi: $2 = $0 + 10
		//           00000000001000100001100000000111
		//mem[2] = 32'b00000000001000100001100000000111; //ADD: $3 = $1 + $2 = 15
		//           01001000000000000000000000000110
		//mem[3] = 32'b01001000000000000000000000000110; //Jal subroutine
		//           
		//mem[4] = 32'b00000100000000000000000000001011; //ADDi: $0 = $0 + 11
		//           00010100011001000000000000000010
		//mem[6] = 32'b00010100011001000000000000000010; //MULi: $4 = $3 * 2 (subroutine)
		//           01001111111000000000000000000000
		//mem[7] = 32'b01001111111000000000000000000000; //JR $ra (bit 31)
		
		
		//*****************--BEQ TEST--******************
		//          000001_00000_00001_0000000000000000
		//mem[0] = 32'b00000100000000010000000000000000;   // ADDi: $1 = $0 + 0
		//          000001_00000_00010_0000000000000001
		//mem[1] = 32'b00000100000000100000000000000001;   // ADDi: $2 = $0 + 1
		//          000001_00000_00011_0000000000001010
		//mem[2] = 32'b00000100000000110000000000000001;   // ADDi: $3 = $0 + 1 (get input)
		//          010100_00011_00010_0000000000000101
		//mem[3] = 32'b01010000011000100000000000001001;   // BEQ: $3 == $2 -> mem[9]
		//	         000001_00000_00001_0000000000001011
		//mem[9] = 32'b00000100000000000000000000001011;   // ADDi: $0 = $0 + 11
		
		//*****************--FIBONACCI--*****************
		//          000001_00000_00000_0000000000000000
		//mem[0] = 32'b00000100000000000000000000000000;   // ADDi: $0 = $0 + 0 //Guarda o valor 0($zero)
		//          000001_00000_00001_0000000000000000
		//mem[1] = 32'b00000100000000010000000000000000;   // ADDi: $1 = $0 + 0 //Guada o F0 = 0
		//          000001_00000_000100000000000000001
		//mem[2] = 32'b00000100000000100000000000000001;   // ADDi: $2 = $0 + 1 //Guarda o F1 = 1
		//          000001_00000_00011_0000000000001010
		//mem[3] = 32'b00000100000000110000000000001010;   // ADDi: $3 = $0 + 10 (TODO: get input)
		//          010100_00011_00000_0000000000001010
		//mem[4] = 32'b01010000011000000000000000001010;   // BEQ: $3 == $0 -> mem[10] --> LOOP Control
		//          000000_00001_00010_00100_00000000000;
		//mem[5] = 32'b00000000001000100010000000000000;   // ADD: $4 = $1 + $2
		//				000000_00010_00000_00001_00000000000
		//mem[6] = 32'b00000000010000000000100000000000;   // ADD: $1 = $2 + $0
		//				000000_00100_00000_00010_00000000000
		//mem[7] = 32'b00000000100000000001000000000000;   // ADD: $2 = $4 + $0
		//				000011_00011_00011_0000000000000001;
		//mem[8] = 32'b00001100011000110000000000000001;   // SUB: $3 = $3 - 1
		//				010001_00000000000000000000000011
		//mem[9] = 32'b01000100000000000000000000000100;   // JUMP: Addr == 4
		//				000001_00000_00000_0000000000001011
		//mem[10]= 32'b00000100000000000000000000001011;   // ADDi: $0 = $0 + 11
		
		
		//*****************--SW(with input)--*****************
		//mem[0] = {16'b0000010000000001, Input[15:0]};      // ADDi: $1 = $0 + 1
		//mem[1] = 32'b100000_00001_00001_0000000000000000;  // SW: $t1, 0($a1)
		//           100000_00001_00001_0000000000000000

		//mem[2] = 32'b011111_00001_00010_0000000000000000;  // LW: $t2, 0($a1)
		//           011111_00001_00010_0000000000000000
