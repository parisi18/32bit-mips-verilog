/*Módulo principal do MIPS 32 bits*/
/*
INSTRUÇÕES SELECIONADAS:
Lógicas:
    - ADD
    - SUB
    - MULT
    - DIV
Aritméticas:
    - AND
    - OR
    - Shift Left
    - Shift Right
Transferência de Dados:
    - LOAD
    - STORE
Branchs condicionais:
    - BEQ
    - BNE
Comparação:
    - SLT
Jump incondicional:
    - JUMP
    - JAL
*/

module ProcessUnit(clk);

input clk;



endmodule