module Registers(clk, rs, rt, rd1, rd2);

input clk;

//
input [4:0] rs, rt;

//Read data 1 e 2
output [31:0] rd1, rd2;

reg [31:0] regs [31:0];



endmodule