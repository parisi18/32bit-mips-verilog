module ALU32(
	input [31:0] a,
	input [31:0] b,
	output [31:0] c
	input [5:0] aluop
);

always(*) begin
	
end

endmodule
