module MemoriaDeInstrucao(addr, inst);

    input [31:0] addr;


endmodule