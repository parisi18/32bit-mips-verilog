module RegisterFile(clk, rs, rt, rd);

input [4:0] rs, rt, rd; 


reg 



endmodule