/*MIPS 32 Instruction Fetching*/

module Pc();



endmodule